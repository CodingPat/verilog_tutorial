module ripple_carry_counter(q,clk,reset);
	output [3:0] q;
	input clk,reset;



